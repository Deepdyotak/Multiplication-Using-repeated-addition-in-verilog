`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.08.2025 20:05:53
// Design Name: 
// Module Name: controlpath
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module controlpath(input clk,eqz,start,
output reg  lda,ldp,clrp,ldb,decb,done);
reg[2:0] state;
parameter S0 = 3'b000, S1 = 3'b001, S2 = 3'b010, S3= 3'b011, S4 = 3'b100;
always@(posedge(clk))begin
case(state)
S0: if(start) state <= S1;
S1: state <= S2;
S2: state<= S3;
S3: #2 if(eqz) state<=S4;
S4: state<=S4;
default: state <= S0;
endcase
end
always@(state) begin
case(state)
S0: begin  #1 lda=0;ldb=0;ldp=0;clrp=0;decb=0; end
S1: begin #1 lda=1; end
S2: begin #1 lda =0; ldb=1; clrp=1; end
S3: begin #1 ldp=1; ldb=0; clrp=0; decb=1; end
S4: begin #1 done=1;ldb=0;ldp=0;decb=0;end
default:begin #1 lda=0;ldb=0;ldp=0;clrp=0;decb=0;end
endcase
end
endmodule
